package axilite_header_pkg ;
  
  `include"../../tb/common/axilite_params.svh"
  
endpackage : axilite_header_pkg