package axilite_scoreboard_pkg;

  // Import all the required packages
  import axilite_trnx_pkg ::* ;
  import axilite_header_pkg ::* ;
  `include"../../tb/scoreboard/axilite_reg_bank.svh"
  `include"../../tb/scoreboard/axilite_comparator.svh"
  `include"../../tb/scoreboard/axilite_predictor.svh"
  `include"../../tb/scoreboard/axilite_scoreboard.svh"

endpackage : axilite_scoreboard_pkg