package axilite_trnx_pkg;
  import axilite_header_pkg :: * ;
  //`include"../../tb/common/axilite_params.svh"
  `include"../../tb/common/transactions/axilite_trnx.svh"

endpackage