package axilite_tx_agent_pkg;

  // Import all the required packages
  import axilite_trnx_pkg ::* ;
  import axilite_header_pkg ::* ;
  

  `include"../../tb/tx_agent/axilite_tx_agt_config.svh"
  `include"../../tb/tx_agent/axilite_generator.svh"
  `include"../../tb/tx_agent/axilite_driver.svh"
  `include"../../tb/tx_agent/axilite_tx_monitor.svh"
  `include"../../tb/tx_agent/axilite_tx_agent.svh"

endpackage