parameter ADDR_WIDTH = 32;
parameter DATA_WIDTH = 32;
parameter logic [31:0] BASEADDR = 32'hA0000000;